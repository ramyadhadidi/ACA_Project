library verilog;
use verilog.vl_types.all;
entity \multiplier__tb\ is
    generic(
        no_of_tests     : integer := 10000
    );
end \multiplier__tb\;
