library verilog;
use verilog.vl_types.all;
entity multiplie_cycle_mips is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
end multiplie_cycle_mips;
