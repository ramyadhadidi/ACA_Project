library verilog;
use verilog.vl_types.all;
entity \single_cycle_mips__tb\ is
    generic(
        end_pc          : integer := 124
    );
end \single_cycle_mips__tb\;
