library verilog;
use verilog.vl_types.all;
entity \multi_cycle_mips__tb\ is
    generic(
        end_pc          : integer := 48
    );
end \multi_cycle_mips__tb\;
