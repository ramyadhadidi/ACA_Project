library verilog;
use verilog.vl_types.all;
entity \pipeline_mips__tb\ is
    generic(
        end_pc          : integer := 48
    );
end \pipeline_mips__tb\;
