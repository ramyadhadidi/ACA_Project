
`timescale 1ns/1ns

module multi_cycle_mips__tb;

	reg clk = 1;
	reg [31:0] counter;
	always @(clk)
		clk <= #5 ~clk;

	reg reset;
	initial begin
		reset = 1;
		counter = 0;
		@(posedge clk);
		@(posedge clk);
		@(posedge clk);
		#1;
		reset = 0;
	end

	initial
		$readmemh("isort32m2.hex", uut.mem.mem_data);

	parameter end_pc = 32'h30;

	integer i;
	always @(uut.pc) begin
	  //$display("counter = %x", counter);
	  counter=counter+1;
		if(uut.pc == end_pc || uut.pc == 32'h20) begin
			for(i=0; i<96; i=i+1) begin
				$write("%x ", uut.mem.mem_data[12+i]);
				if(((i+1) % 16) == 0)
					$write("\n");
			end
			$stop;
		end
	end

	multi_cycle_mips uut(
		.clk(clk),
		.reset(reset)
	);


endmodule

