library verilog;
use verilog.vl_types.all;
entity async_mem is
    port(
        clk             : in     vl_logic;
        write           : in     vl_logic;
        address         : in     vl_logic_vector(31 downto 0);
        write_data      : in     vl_logic_vector(31 downto 0);
        read_data       : out    vl_logic_vector(31 downto 0)
    );
end async_mem;
